LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY alu_tb IS
END alu_tb;

ARCHITECTURE alu_tb_arch OF alu_tb IS

CONSTANT N_USER: INTEGER := 4;

COMPONENT alu
	GENERIC(N: INTEGER := 4);
	PORT(A_BUS, B_BUS: IN SIGNED(N-1 DOWNTO 0); 					--Inputs
		  F_BUS: IN STD_LOGIC_VECTOR(2 DOWNTO 0);			 		--Select
		  CBin: IN STD_LOGIC;									 		--Carry/Borrow In
		  C_BUS: OUT SIGNED(N-1 DOWNTO 0);		 					--Output
		  CBout: OUT STD_LOGIC;								    		--Carry/Borrow Out
		  A_SSD, B_SSD, C_SSD: OUT STD_LOGIC_VECTOR(0 TO 6);	--Hex Decimal Displays
		  A_NEG, B_NEG, C_NEG: OUT STD_LOGIC_VECTOR(0 TO 6);	--Hex Negative Displays
		  OV_SEG: OUT STD_LOGIC_VECTOR(0 TO 6);					--Hex Overflow Display
		  CBout_SEG: OUT STD_LOGIC_VECTOR(0 TO 6);				--Hex Carry/Borrow Out
		  CBin_LED: OUT STD_LOGIC;										--LED Carry/Borrow In
		  OVERFLOW: OUT STD_LOGIC);									--Overflow
END COMPONENT;

SIGNAL ABUSTEST, BBUSTEST, CBUSTEST: SIGNED(N_USER-1 DOWNTO 0);
SIGNAL CBINTEST, CBOUTTEST, OVTEST: STD_LOGIC;
SIGNAL FBUSTEST: STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN
U1: alu PORT MAP (ABUSTEST, BBUSTEST, FBUSTEST, CBINTEST, CBUSTEST, CBOUTTEST, OVERFLOW => OVTEST); 

ABUSTEST <= "0110";
BBUSTEST <= "0011";
CBINTEST <= '1';

PROCESS
	BEGIN
		FBUSTEST <= "000";
		WAIT FOR 20ns;
		FBUSTEST <= "001";
		WAIT FOR 20ns;
		FBUSTEST <= "010";
		WAIT FOR 20ns;
		FBUSTEST <= "011";
		WAIT FOR 20ns;
		FBUSTEST <= "100";
		WAIT FOR 20ns;
		FBUSTEST <= "101";
		WAIT FOR 20ns;
		FBUSTEST <= "110";
		WAIT FOR 20ns;
		FBUSTEST <= "111";
		WAIT FOR 20ns;
END PROCESS; 
  
END alu_tb_arch;

