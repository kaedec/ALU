LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RCA_4bit IS

	PORT(A, B: IN SIGNED(3 DOWNTO 0);
			C0: IN STD_LOGIC;
			S: OUT SIGNED(3 DOWNTO 0);
			C4, OV: OUT STD_LOGIC);
END RCA_4bit;

ARCHITECTURE RCA_4bit_arch OF RCA_4bit IS

COMPONENT and_gate PORT (A, B: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT inverter PORT(A: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT or_gate PORT(A, B: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT xor_struct PORT (A, B: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT xor_gate_3i PORT (A, B, C: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT or_gate_3i PORT (A, B, C: IN STD_LOGIC; F: OUT STD_LOGIC);
	END COMPONENT;
	
COMPONENT full_adder PORT (A, B, Cin: IN STD_LOGIC; Sum, Cout: OUT STD_LOGIC);
	END COMPONENT;
	
SIGNAL C1, C2, C3, C4_ov: STD_LOGIC;

BEGIN

U1: full_adder PORT MAP(A(0), B(0), C0, S(0), C1);
U2: full_adder PORT MAP(A(1), B(1), C1, s(1), C2);
U3: full_adder PORT MAP(A(2), B(2), C2, s(2), C3);
U4: full_adder PORT MAP(A(3), B(3), C3, s(3), C4_ov);
U5: xor_struct PORT MAP(C3, C4_ov, OV);

C4 <= C4_ov;

END RCA_4bit_arch;